attribute ASYNC_REG : string;
attribute ASYNC_REG of sync_regs: signal is "TRUE";