attribute fsm_encoding : string;
attribute fsm_encoding of state : signal is "gray";
