constant rom : ram_type;