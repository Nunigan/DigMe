constant constant_name : type := value; -- Definition
constant countersize : integer := 2**16-1; -- Example 1
constant cmdreadid : std_logic_vector(7 downto 0) := x"9F"; -- Example 2