attribute ram_style : string;
attribute ram_style of blockram : variable is "block";