constant ROM : rom_type :=("00000000", "00000011", ..., "00100000")