attribute fsm_safe_state : string;
attribute fsm_safe_state of state : signal is "reset_state";
