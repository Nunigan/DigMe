attribute keep_hierarchy : string;
attribute keep_hierarchy of beh : architecture is "yes";