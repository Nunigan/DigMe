use work.my_package.all;